/* *********************************************
This file is a top module to generate clk, rst and start signal
************************************************ */


module clk_rst();

reg clk;
reg rst;
reg start;
reg halt;


always begin
    clk <= 'd0;
    #1;
    clk <= ~clk;
    #1;
end

initial begin
    rst <= 'd1;
    start <= 'd0;
    halt <= 'd0;
    #5;
    rst <= 'd0;
    #2;
    start <= 'd1;
    #2;
    start <= 'd0;
    #2;
    #2;
    #2;
    // halt <= 'd1;
    // #2;
    // halt <= 'd0;
end


// initial begin
//     rst <= 'd1;
//     start <= 'd0;
//     need_data <= 'd0;
//     #5;
//     rst <= 'd0;
//     #2;
//     start <= 'd1;
//     #2;
//     start <= 'd0;
//     #2;
//     need_data <= 'd1;
//     #2;
//     need_data <= 'd0;
//     #20;
//     need_data <= 'd1;
//     #2;
//     need_data <= 'd0;
// end

CONV1_LAYER1_DENSE_TOP conv1_layer1_dense_top(
    .clk                        (clk),
    .rst                        (rst),
    .start                      (start),
    .halt                       (halt)
);


// wire                                                reg_data_v_w;
// wire    [1023:0]                                    reg_data_w;
// reg                                                 data_v;
// reg     [1023:0]                                    in_veca_data;
// reg     [15:0]                                      in_sig_data;
// reg                                                 usr_rst;


// initial begin
//     rst <= 'd1;
//     data_v <= 'd0;
//     usr_rst <= 'd0;
//     #5;
//     rst <= 'd0;
//     #2;
//     data_v <= 'd1;
//     #2;
//     data_v <= 'd1;
//     #2;
//     data_v <= 'd1;
//     #2;
//     data_v <= 'd1;
//     #2;
//     data_v <= 'd1;
//     #2;
//     data_v <= 'd1;
//     #2;
//     data_v <= 'd0;

//     #200;
//     usr_rst <= 'd1;
    
//     #2;
//     data_v <= 'd1;
//     usr_rst <= 'd0;
//     #2;
//     data_v <= 'd0;
//     #2;
// end

// always @ (posedge clk) begin
//     in_sig_data <= 'h0100;
//     in_veca_data <= 'h0100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100010001000100;
// end


// TB4PARAMULT_REGHEAP tb4paramult_regheap(
//     .clk                                (clk),
//     .rst                                (rst),
//     .data_v                             (data_v),
//     .in_veca_data                       (in_veca_data),
//     .in_sig_data                        (in_sig_data),
//     .usr_rst                            (usr_rst),
//     .reg_data_w                         (reg_data_w),
//     .reg_data_v_w                       (reg_data_v_w)
// );




// reg     [95:0]                          in_fea;
// reg     [95:0]                          in_wei;
// reg     [5:0]                           non_zero;


// initial begin
//     rst <= 'd1;
//     #2;
//     rst <= 'd0;
//     #10;
//     in_fea <= 96'h0600_0500_0400_0300_0200_0100;
//     in_wei <= 96'h0600_0500_0400_0300_0200_0100;
//     // non_zero <= 6'b111_111;
//     // #2;
//     non_zero <= 6'b111_010;
//     #2;
//     non_zero <= 6'b001_111;
//     #2;
//     non_zero <= 6'b101_101;
//     #2;
//     // non_zero <= 6'b000_000;
//     // #2;
//     non_zero <= 6'b000_000;

// end







// DYN_ISSUE demo(
//     .clk                                (clk),
//     .rst                                (rst),
//     .in_fea                             (in_fea),
//     .in_wei                             (in_wei),
//     .non_zero                           (non_zero)
// );


endmodule



